// add 3, 1-bits
module FAdder(output reg carry, sum, input a, b, c);
  always @ (*) begin
    
  end  
