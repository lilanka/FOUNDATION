module KY32_imem(
  output  [31:0]  ins,
  input   [31:0]  a
);

  wire  [31:0]  imem [0:31] // 1MB
endmodule
