`include "ram.v"

module Memory(out, in, addr, clk, ld);
  input [15:0] in;
  input [14:0]
  

Economic 




















































